
module expand(z,x,y);
input x,y;
output z;
and a_1(z,x,y);
end module